package max_tb_tasks;





endpackage